// ******************************************************************
// Specific defines needed for building
// ******************************************************************

`define WT_DCACHE // use the write-through cache by default
`define DISABLE_TRACER // remove the default tracer widget
`define SRAM_NO_INIT // disable setting srams
